`include "mycpu.h"

module exe_stage(
    input                          clk           ,
    input                          reset         ,
    //allowin
    input                          ms_allowin    ,
    output                         es_allowin    ,
    //from ds
    input                          ds_to_es_valid,
    input  [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus  ,
    //to ms
    output                         es_to_ms_valid,
    output [`ES_TO_MS_BUS_WD -1:0] es_to_ms_bus  ,
    // data sram interface
    output        data_sram_en   ,
    output [ 3:0] data_sram_wen  ,
    output [31:0] data_sram_addr ,
    output [31:0] data_sram_wdata,
    output [ 4:0] es_real_dest,
    output [31:0] exe_forward_data,
    output        es_res_from_mem,
    output [31:0] exe_forward_data_HI,//lab6
    output [31:0] exe_forward_data_LO,//lab6
    output        es_mt_op,
    output        es_mult_multu_div_divu_op,
    output [`SPECIAL_REG_ADDR_WD -1:0] es_dest_special
);

reg         es_valid      ;
wire        es_ready_go   ;

reg  [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus_r;
wire [15:0] es_alu_op     ;
wire        es_load_op    ;
wire        es_mf_op      ;//lab6
//wire        es_mt_op      ;//lab6
//wire        es_mult_multu_div_divu_op;//lab6
wire        es_src1_is_sa ;  
wire        es_src1_is_pc ;
wire        es_src2_is_imm_signextend;
wire        es_src2_is_imm_zeroextend;
wire        es_src2_is_8  ;
wire        es_gr_we      ;
wire        es_mem_we     ;
wire [ 4:0] es_dest       ;
//wire [`SPECIAL_REG_ADDR_WD -1:0] es_dest_special;//lab6
wire [15:0] es_imm        ;
wire [31:0] es_rs_value   ;
wire [31:0] es_rt_value   ;
wire [31:0] es_special_value;//lab6
wire [31:0] es_pc         ;
assign {
        es_mult_multu_div_divu_op   ,  //177:177 lab6
        es_mt_op                    ,  //176:176 lab6
        es_special_value            ,  //175:144 lab6
        es_mf_op                    ,  //143:143 lab6
        es_dest_special             ,  //142:141 lab6
        es_src2_is_imm_zeroextend   ,  //140:140
        es_alu_op                   ,  //139:124
        es_load_op                  ,  //123:123
        es_src1_is_sa               ,  //122:122
        es_src1_is_pc               ,  //121:121
        es_src2_is_imm_signextend   ,  //120:120
        es_src2_is_8                ,  //119:119
        es_gr_we                    ,  //118:118
        es_mem_we                   ,  //117:117
        es_dest                     ,  //116:112
        es_imm                      ,  //111:96
        es_rs_value                 ,  //95 :64
        es_rt_value                 ,  //63 :32
        es_pc                          //31 :0
       } = ds_to_es_bus_r;

wire [31:0] es_alu_src1   ;
wire [31:0] es_alu_src2   ;
wire [31:0] es_alu_result ;
wire [31:0] es_alu_result_HI;//lab6

wire    unsigned_dout_tvalid;
wire    signed_dout_tvalid;  

//wire        es_res_from_mem;//lab5 changed
wire        es_res_from_special;//lab6
wire        es_res_from_rs;//lab6

assign es_res_from_mem = es_load_op;
assign es_res_from_special = es_mf_op;//lab6
assign es_res_from_rs = es_mt_op;//lab6
assign es_to_ms_bus = {
                        es_mult_multu_div_divu_op, //171:171 lab6
                        es_rs_value             ,  //170:139 lab6
                        es_res_from_rs          ,  //138:138 lab6
                        es_alu_result_HI        ,  //137:106 lab6
                        es_special_value        ,  //105:74 lab6
                        es_res_from_special     ,  //73:73 lab6
                        es_dest_special         ,  //72:71 lab6
                        es_res_from_mem         ,  //70:70
                        es_gr_we                ,  //69:69
                        es_dest                 ,  //68:64
                        es_alu_result           ,  //63:32
                        es_pc                      //31:0
                        };

//assign es_ready_go    = (alu_op[14]) ? !signed_dout_tvalid  : 1'b1;
assign es_ready_go    = ~((es_alu_op[14] && !signed_dout_tvalid) || (es_alu_op[15] && !unsigned_dout_tvalid));



assign es_allowin     = !es_valid || es_ready_go && ms_allowin;
assign es_to_ms_valid =  es_valid && es_ready_go;
always @(posedge clk) begin
    if (reset) begin
        es_valid <= 1'b0;
    end
    else if (es_allowin) begin
        es_valid <= ds_to_es_valid;
    end

    if (ds_to_es_valid && es_allowin) begin
        ds_to_es_bus_r <= ds_to_es_bus;
    end
end

assign es_alu_src1 = es_src1_is_sa  ? {27'b0, es_imm[10:6]} : 
                     es_src1_is_pc  ? es_pc[31:0] :
                                      es_rs_value;
assign es_alu_src2 =
                    es_src2_is_imm_signextend ? {{16{es_imm[15]}}, es_imm[15:0]} :
                    es_src2_is_imm_zeroextend ? {{16{1'b0}}, es_imm[15:0]} ://lab6 new
                    es_src2_is_8   ? 32'd8 :
                    es_rt_value;

alu u_alu(
    .clk        (clk),
    .reset      (reset),
    .signed_dout_tvalid (signed_dout_tvalid),
    .unsigned_dout_tvalid   (unsigned_dout_tvalid),
    .alu_op     (es_alu_op    ),
    .alu_src1   (es_alu_src1  ),
    .alu_src2   (es_alu_src2  ),
    .alu_result (es_alu_result),
    .alu_result_HI (es_alu_result_HI)//lab6
    );

assign data_sram_en    = 1'b1;
assign data_sram_wen   = es_mem_we&&es_valid ? 4'hf : 4'h0;
assign data_sram_addr  = es_alu_result;
assign data_sram_wdata = es_rt_value;
assign es_real_dest = (es_valid & es_gr_we) ? es_dest : 5'b00000;//if no inst, let real_dest be 0.
assign exe_forward_data = es_alu_result;//lab5
assign exe_forward_data_HI = es_mt_op ? es_rs_value : es_alu_result_HI;//lab6
assign exe_forward_data_LO = es_mt_op ? es_rs_value : es_alu_result;//lab6

endmodule